// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	CoinsMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input	logic	[10:0] offsetX,// offset from top left  position 
					input	logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket
					input	logic	coinCollision,
					input logic [4:0] randomMapLocationX,
					input logic [3:0] randomMapLocationY,
					input logic placeCoin,		// a pulse evrey 2 sec
					input logic placeMoneyBag,	// a pulse evrey 4 sec
					input logic placeTimeBoost,	// a pulse evrey 20 sec

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
					output	logic upScore,			// pulse when pacman eats money bag
					output	logic upTime			// pulse when pacman eats time boost
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel
localparam  int MAZE_NUMBER_OF_X_LOGICS = 18;
localparam  int MAZE_NUMBER_OF_Y_LOGICS = 12;     


// flags that are in charge of looking for a different spot to place coins and money bags
logic pick_anotherCoin_flag ; // goes up if the spot for the coin is already taken
logic pick_anotherMoneyBag_flag ;


// if the random map Y location is greater than 11, take only the 3 lower bits
logic [3:0] Y_adjustment ;
assign Y_adjustment = (randomMapLocationY[3] & randomMapLocationY[2]) ? {1'b0,randomMapLocationY[2:0]} : randomMapLocationY[3:0] ;


// the playing screen is 576*384  or  18 * 12 squares of 32*32  bits 
logic [0:MAZE_NUMBER_OF_Y_LOGICS-1] [0:MAZE_NUMBER_OF_X_LOGICS-1] [2:0] MazeBitMapMask ;


// specifies the starting value needed for each square
// this bit map will load to the playing bit map on evrey reset
// 3'h004 marks a place where no wall could be placed

/* FOR TESTING */
/*
logic [0:MAZE_NUMBER_OF_Y_LOGICS-1] [0:MAZE_NUMBER_OF_X_LOGICS-1] [2:0]  starting_MazeBitMapMask= 
{{3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00},
 {3'h00, 3'h04, 3'h04, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00},
 {3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00},
 {3'h04, 3'h04, 3'h04, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h04, 3'h04},
 {3'h00, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h00},
 {3'h00, 3'h04, 3'h00, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h04, 3'h03, 3'h04, 3'h00},
 {3'h00, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h04, 3'h00},
 {3'h00, 3'h04, 3'h00, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00},
 {3'h00, 3'h04, 3'h00, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00},
 {3'h00, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00},
 {3'h00, 3'h04, 3'h00, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00, 3'h00, 3'h04, 3'h04, 3'h00},
 {3'h00, 3'h00, 3'h00, 3'h04, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00, 3'h00}
 };
*/

logic [0:MAZE_NUMBER_OF_Y_LOGICS-1] [0:MAZE_NUMBER_OF_X_LOGICS-1] [2:0]  starting_MazeBitMapMask= 
{{3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01},
 {3'h01, 3'h04, 3'h04, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h04, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01},
 {3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01},
 {3'h04, 3'h04, 3'h04, 3'h04, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h04, 3'h04, 3'h04, 3'h04},
 {3'h02, 3'h02, 3'h02, 3'h04, 3'h01, 3'h01, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h04, 3'h01, 3'h01, 3'h04, 3'h01, 3'h01, 3'h01},
 {3'h02, 3'h04, 3'h02, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h04, 3'h01, 3'h04, 3'h01},
 {3'h02, 3'h02, 3'h02, 3'h04, 3'h01, 3'h01, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h04, 3'h01, 3'h01, 3'h04, 3'h04, 3'h04, 3'h01},
 {3'h02, 3'h04, 3'h02, 3'h04, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01},
 {3'h02, 3'h04, 3'h02, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01},
 {3'h02, 3'h02, 3'h02, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01},
 {3'h02, 3'h04, 3'h02, 3'h01, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01, 3'h01, 3'h04, 3'h04, 3'h01},
 {3'h02, 3'h02, 3'h02, 3'h04, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01, 3'h01}
 };


 logic [0:2] [0:31] [0:31] [7:0]  object_colors  = {
 // coins bitmap
{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hf8,8'hf8,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hf8,8'hfd,8'hfd,8'hf8,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hf8,8'hfd,8'hf9,8'hf8,8'hf9,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf9,8'hf8,8'hf8,8'hf8,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf9,8'hf9,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
},

// money bag
{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6c,8'h8c,8'h8c,8'hd9,8'hf9,8'hf9,8'hd9,8'hf8,8'h8d,8'h8c,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf9,8'hf9,8'hfe,8'hd4,8'hb4,8'hd4,8'hb4,8'hd4,8'hfe,8'hfd,8'hf9,8'h6c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'h00,8'hb4,8'h90,8'h90,8'h90,8'hd5,8'h00,8'hb4,8'hf9,8'h6c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf9,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf9,8'hf9,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd9,8'hd4,8'hd9,8'hf9,8'hf9,8'hf9,8'hf9,8'hb4,8'hd9,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6c,8'h90,8'hf9,8'hf9,8'hb4,8'h00,8'hd4,8'h90,8'hd4,8'hd4,8'hf9,8'h90,8'hd5,8'h00,8'hb4,8'hf9,8'hf9,8'hf9,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf9,8'hd8,8'hd4,8'hd4,8'hb4,8'h90,8'h00,8'h00,8'h90,8'hd9,8'hb0,8'h00,8'h00,8'hd5,8'hfd,8'hf9,8'hf9,8'hfe,8'hd9,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hd4,8'hd4,8'hb4,8'hb4,8'h90,8'hd4,8'h90,8'h90,8'h00,8'h00,8'h00,8'h90,8'h90,8'hfd,8'hfe,8'hfe,8'hfe,8'hd9,8'hfe,8'hf9,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hd4,8'hd4,8'hb4,8'h8c,8'hd4,8'hd4,8'hf9,8'hd4,8'h90,8'hb0,8'h8c,8'hf9,8'hf9,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hf9,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'hd4,8'hb0,8'h8c,8'hd4,8'hd4,8'hd4,8'hb4,8'hf9,8'h00,8'hd9,8'h00,8'hf9,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hf9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'h90,8'hb0,8'hd4,8'h8c,8'hb4,8'hd4,8'hf9,8'hd4,8'h00,8'hfd,8'h00,8'hf9,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hf9,8'hfe,8'hfd,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'hb4,8'hd9,8'hb4,8'hd4,8'hb4,8'hd4,8'hb4,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hf9,8'hd9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'h90,8'hd9,8'hf9,8'hb4,8'hb0,8'hb4,8'h00,8'hd4,8'h00,8'hd9,8'h00,8'hfe,8'h00,8'hfe,8'hfe,8'hfa,8'hfd,8'hfe,8'hd9,8'hfd,8'hd9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'hd4,8'hb0,8'h90,8'hb4,8'h90,8'hd4,8'h00,8'hd9,8'h00,8'hd9,8'h00,8'hfe,8'h00,8'hfe,8'hf9,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'hb0,8'hb4,8'hd4,8'h8c,8'hd4,8'hd4,8'hd4,8'h00,8'h00,8'hb4,8'h00,8'hd9,8'hf9,8'hf9,8'hf9,8'hf9,8'hfd,8'hd9,8'hd9,8'hd9,8'hf9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'hd4,8'hb4,8'h90,8'hd4,8'h90,8'hd4,8'hd4,8'hb4,8'h00,8'h00,8'h00,8'hd9,8'hf9,8'hd9,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hd4,8'hf9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'h90,8'hb0,8'hd4,8'h90,8'hd4,8'h90,8'hb4,8'hb4,8'h00,8'hd4,8'h00,8'h00,8'hd9,8'hb4,8'hf9,8'hd4,8'hd4,8'hf9,8'hd4,8'hf9,8'hd9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'hd4,8'hb0,8'h90,8'hd4,8'h90,8'hd4,8'h00,8'hd4,8'h00,8'hd4,8'h00,8'hd9,8'h00,8'hf9,8'hb4,8'hf9,8'hf9,8'hd4,8'hd9,8'hd4,8'hd9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'hd9,8'hb4,8'hd4,8'hd4,8'hb4,8'h8c,8'hd4,8'h90,8'h00,8'h90,8'h00,8'hb4,8'h00,8'hb4,8'h00,8'hd5,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd9,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'h24,8'h8c,8'hd4,8'hb4,8'h8c,8'hd4,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb4,8'hb4,8'hb4,8'hd4,8'hd0,8'hb4,8'h00,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'hd5,8'h90,8'h24,8'h00,8'hd4,8'hb4,8'h90,8'hd4,8'h90,8'h00,8'h90,8'h00,8'h90,8'hd4,8'hb0,8'hd4,8'hd4,8'hd5,8'h00,8'hb0,8'hb4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'h24,8'h8c,8'hd4,8'h90,8'h90,8'hd4,8'h90,8'hb4,8'h00,8'hd4,8'h00,8'hb0,8'hb0,8'hd4,8'h90,8'h90,8'h90,8'hb4,8'h00,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd5,8'hb4,8'hd4,8'hd4,8'hb4,8'h90,8'h90,8'h90,8'h90,8'h90,8'h90,8'hb0,8'h90,8'h90,8'hd4,8'hd4,8'hb0,8'hd4,8'hb4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
},

// time boost
{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h64,8'h6c,8'h6c,8'h64,8'h64,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hcc,8'hf8,8'hf8,8'hfc,8'hfc,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h64,8'hf0,8'hd0,8'h24,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6c,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h60,8'ha0,8'ha0,8'ha0,8'ha0,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h60,8'h80,8'ha0,8'ha4,8'hd6,8'hd6,8'ha0,8'hc0,8'h80,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h60,8'ha0,8'hac,8'hfa,8'hff,8'hff,8'h00,8'hff,8'hd1,8'ha4,8'hc0,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hd1,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'had,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'ha4,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hd6,8'hc0,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'ha0,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'ha4,8'hc0,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h80,8'hff,8'h00,8'hff,8'hff,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'h00,8'hfa,8'ha0,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h80,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'ha4,8'ha0,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'ha0,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'ha4,8'ha0,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'ha0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hd6,8'hc0,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hd1,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h60,8'ha0,8'ha4,8'hfa,8'hff,8'h00,8'h00,8'hff,8'hd5,8'ha4,8'hc0,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h60,8'h80,8'ha0,8'h84,8'hd1,8'hd1,8'ha0,8'hc0,8'h80,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h60,8'ha0,8'ha0,8'ha0,8'ha0,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
}};
 
//////////--------------------------------------------------------------------------------------------------------------= 

// pipeline (ff) to get the pixel color from the array 	 

//----------------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask <= starting_MazeBitMapMask ;
	end // resetN
	
	else begin
		// defaults
		RGBout <= TRANSPARENT_ENCODING ; 
		MazeBitMapMask <= MazeBitMapMask ;
		pick_anotherCoin_flag <= 1'b0 ;
		pick_anotherMoneyBag_flag <= 1'b0 ; 
		upScore <= 1'b0 ;
		upTime <= 1'b0 ;
		// end of defaults
		
		// coins drawing and deleting
		if (InsideRectangle == 1'b1 ) begin
			case (MazeBitMapMask[offsetY[8:5]][offsetX[9:5]])
				3'h01 : RGBout <= object_colors [0][offsetY[4:0]][offsetX[4:0]] ;	// regular coin
				3'h02 : RGBout <= object_colors [1][offsetY[4:0]][offsetX[4:0]] ;	// money bag
				3'h03 : RGBout <= object_colors [2][offsetY[4:0]][offsetX[4:0]] ;	// time boost
				default: RGBout <= TRANSPARENT_ENCODING ;
			endcase


				
			if (coinCollision == 1'b1) begin									 // if pacman touches a coin
				MazeBitMapMask[offsetY[8:5]][offsetX[9:5]] <= 0	;		// the coin will stop showing
				case (MazeBitMapMask[offsetY[8:5]][offsetX[9:5]])
					3'h02 : upScore <= 1'b1 ;
					3'h03 : upTime <= 1'b1 ;
					default: begin
									upScore <= 1'b0 ;
									upTime <= 1'b0 ;
					end // default
				endcase
			end
		end // InsideRectangle
		
		
		// set the conditions to add a coins to the game
		// regular coins logic
		if ( placeCoin	|| pick_anotherCoin_flag ) begin	
			if (MazeBitMapMask[Y_adjustment[3:0]][randomMapLocationX[4:0]] == 0) begin
				MazeBitMapMask[Y_adjustment[3:0]][randomMapLocationX[4:0]] <= 3'h01;
				pick_anotherCoin_flag <= 1'b0 ;
			end
			else pick_anotherCoin_flag <= 1'b1;
		end // placeCoin || pick_anotherCoins_flag

		
		// money bags logic
		if ( placeMoneyBag	|| pick_anotherMoneyBag_flag ) begin	
			if (MazeBitMapMask[Y_adjustment[3:0]][randomMapLocationX[4:0]] == 0) begin
				MazeBitMapMask[Y_adjustment[3:0]][randomMapLocationX[4:0]] <= 3'h02;
				pick_anotherMoneyBag_flag <= 1'b0;
			end
			else pick_anotherMoneyBag_flag <= 1'b1;
					
		end // placeMoneyBag || pick_anotherMoneyBag_flag
		
		
		// time boost logic
		if ( placeTimeBoost == 1'b1 )
			MazeBitMapMask[5][15] <= 4'h03;
	 
	end // else statement
end // always_ff

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

